*Obem_Att_1dB
Vg 1 0 AC 1

Rg 1 25 0.01

*RA12 27 0 465.2
*RA13 27 7 930.4
*RA14 27 2 476

RB21 25 2 1.44
RB23 2 8 2.88
RB24 2 3 2.88


RC31 25 3 1.44
RC33 3 9 2.88
RC34 3 4 2.88

RD41 25 4 1.44
RD43 4 10 2.88
RD44 4 5 2.88

RE51 25 5 1.44
RE53 5 11 2.88
RE54 5 6 435.4

RF63 6 12 868
RF64 6 0 434

*RG12 7 0 465.2
*RG13 7 13 930.4
*RG14 7 8 476.5

RH23 8 14 2.88
RH24 8 9 2.88

RL33 9 15 2.88
RL34 9 10 2.88

RM43 10 16 2.88
RM44 10 11 2288

RN53 11 17 2.88
RN54 11 12 435.4

RO63 12 18 868
RO64 12 0 434

*RP12 13 0 465.2
*RP13 13 19 930.4
*RP14 13 14 476.5

RR23 14 20 2.88
RR24 14 15 2.88

RS33 15 21 2.88
RS34 15 16 2.88

RJ43 16 22 2.88
RJ44 16 17 2.88

RK53 17 23 2.88
RK54 17 18 435.4

RV63 18 24 868
RV64 18 0 434

*RI12 19 0 465.2
*RI14 19 20 476.5

RQ23 20 26 1.44
RQ24 20 21 2.88

RW33  21 26 1.44
RW34 21 22 2.88

RT43 22 26 1.44
RT44 22 23 2.88

RY53 23 26 1.44
RY54 23 24 435.4

RZ64 24 0 434



Rout 26 0 50



.PROBE
*.Tran 0 1 1m
.AC LIN  1000 100 200
*.DC LIN 1000
.END
